
class my_agent extends uvm_agent;


    `uvm_component_utils(my_agent)
    
    my_driver drv;
    my_sequencer seqr;
    
    function new(string name, uvm_component parent);
        super.new(name, parent);
    endfunction
    
    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        seqr = my_sequencer::type_id::create("seqr", this);
        drv = my_driver::type_id::create("drv", this);
    endfunction

    function void connect_phase(uvm_phase phase);
        drv.seq_item_port.connect(seqr.seq_item_export);
    endfunction

endclass